module tank(input logic Reset, GReset, frame_clk, tank,
				input logic [7:0] keycode,
				output logic  [9:0] TankX, TankY, TankSize, TankXMot, TankYMot);
				
	logic [9:0] Tank_X_Pos, Tank_X_Motion, Tank_Y_Pos, Tank_Y_Motion, Tank_Size;
	 
    parameter [9:0] Tank_X_Center=640;  // Center position on the X axis
    parameter [9:0] Tank_Y_Center=480;  // Center position on the Y axis
    parameter [9:0] Tank_X_Min=16;       // Leftmost point on the X axis
    parameter [9:0] Tank_X_Max=623;     // Rightmost point on the X axis
    parameter [9:0] Tank_Y_Min=55;       // Topmost point on the Y axis
    parameter [9:0] Tank_Y_Max=465;     // Bottommost point on the Y axis
    parameter [9:0] Tank_X_Step=1;      // Step size on the X axis
    parameter [9:0] Tank_Y_Step=1;      // Step size on the Y axis

    assign Tank_Size = 16;  // assigns the value 4 as a 10-digit binary number, ie "0000000100"
   
    always_ff @ (posedge Reset or posedge frame_clk or posedge GReset )
    begin: Move_Ball
        if (Reset)  // Asynchronous Reset
        begin 
            Tank_Y_Motion <= 10'd0; //Ball_Y_Step;
				Tank_X_Motion <= 10'd0; //Ball_X_Step;
				Tank_Y_Pos <= Tank_Y_Center;
				Tank_X_Pos <= Tank_X_Center;
        end
        else if (GReset)
		  begin
				Tank_Y_Motion <= 10'd0; //Ball_Y_Step;
				Tank_X_Motion <= 10'd0; //Ball_X_Step;
				Tank_Y_Pos <= Tank_Y_Center;
				Tank_X_Pos <= Tank_X_Center;
		  end
        else
		  
        begin
		  
				 if ( (Tank_Y_Pos + Tank_Size) >= Tank_Y_Max )  // Ball is at the bottom edge, BOUNCE!
					  Tank_Y_Motion <= 0;  // 2's complement.
					  
				 if ( (Tank_Y_Pos - Tank_Size) <= Tank_Y_Min )  // Tank is at the top edge, BOUNCE!
					  Tank_Y_Motion <= 0;
					  
				 if ( (Tank_X_Pos + Tank_Size) >= Tank_X_Max )  // Tank is at the Right edge, BOUNCE!
					  Tank_X_Motion <= 0;  // 2's complement.
					  
				 if ( (Tank_X_Pos - Tank_Size) <= Tank_X_Min )  // Tank is at the Left edge, BOUNCE!
					  Tank_X_Motion <= 0;
				 case (keycode)
					8'h04 : begin
								if (tank == 0)
								begin
									if (((Tank_X_Pos - Tank_Size) > Tank_X_Min))
									begin
										Tank_X_Motion <= -1;//A
										Tank_Y_Motion<= 0;
									end
								end
							  end
					        
					8'h07 : begin
							  if (tank == 0)
							  begin
									if (~((Tank_X_Pos + Tank_Size)+1 >= Tank_X_Max))
									begin
										Tank_X_Motion <= 1;//D
										Tank_Y_Motion <= 0;
									end
							  end
							  end

							  
					8'h16 : begin
								if (tank == 0)
								begin
									if (~((Tank_Y_Pos + Tank_Size)+1 >= Tank_Y_Max ))
									begin
										Tank_Y_Motion <= 1;//S
										Tank_X_Motion <= 0;
									end
							  end
							 end
							  
					8'h1A : begin
								if (tank == 0)
								begin
									if(((Tank_Y_Pos - Tank_Size) > Tank_Y_Min ))
									begin
									Tank_Y_Motion <= -1;//W
									Tank_X_Motion <= 0;
									end
							  end
							 end
					8'h0d : begin
								if (tank == 1)
								begin
									if (((Tank_X_Pos - Tank_Size) > Tank_X_Min))
									begin
										Tank_X_Motion <= -1;//A
										Tank_Y_Motion<= 0;
									end
								end
							  end
					        
					8'h0f : begin
							  if (tank == 1)
							  begin
								if (~((Tank_X_Pos + Tank_Size)+1 >= Tank_X_Max))
									begin
										Tank_X_Motion <= 1;//D
										Tank_Y_Motion <= 0;
									end
							  end
							  end

							  
					8'h0e : begin
								if (tank == 1)
								begin
									if (~((Tank_Y_Pos + Tank_Size)+1 >= Tank_Y_Max ))
									begin
									Tank_Y_Motion <= 1;//S
									Tank_X_Motion <= 0;
									end
							  end
							 end
							  
					8'h0c : begin
								if (tank == 1)
								begin
									if(((Tank_Y_Pos - Tank_Size) > Tank_Y_Min ))
									begin
										Tank_Y_Motion <= -1;//W
										Tank_X_Motion <= 0;
									end
							  end
							 end		 
					default: ;
			   endcase 	  

					  
				 
				 
				 
				 Tank_Y_Pos <= (Tank_Y_Pos + Tank_Y_Motion);  // Update Tank position
				 Tank_X_Pos <= (Tank_X_Pos + Tank_X_Motion);
			
			
	  /**************************************************************************************
	    ATTENTION! Please answer the following quesiton in your lab report! Points will be allocated for the answers!
		 Hidden Question #2/2:
          Note that Ball_Y_Motion in the above statement may have been changed at the same clock edge
          that is causing the assignment of Ball_Y_pos.  Will the new value of Ball_Y_Motion be used,
          or the old?  How will this impact behavior of the ball during a bounce, and how might that 
          interact with a response to a keypress?  Can you fix it?  Give an answer in your Post-Lab.
      **************************************************************************************/
      
			
		end  
    end
       
    assign TankX = Tank_X_Pos;
   
    assign TankY = Tank_Y_Pos;
   
    assign TankSize = Tank_Size;
    
	 assign TankXMot = Tank_X_Motion;
	 
	 assign TankYMot = Tank_Y_Motion;

endmodule
